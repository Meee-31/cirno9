`include "cirno9_define.v"

module cirno9_core(
    input         rst_n,
    input         clk,
);
endmodule