`include "cirno9_define.v"

module cirno9_core(
    input         rst_n,
    input         clk,
    
    output [31:0] o_itcm_adr,
    input  [31:0] i_intm_dat,
);
endmodule